// Honzales top module
// Copyright 2022 Andreas Wendleder

module honzales();
        initial begin
                $display("honzales starts");
        end
endmodule

